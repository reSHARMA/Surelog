module foo #(localparam happy_lp=1)
  (output o);
  assign o = happy_lp;
endmodule
