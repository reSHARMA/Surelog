module test (input size);
    logic [size:0] foo [size-1 : 0];
endmodule
