module foo (input i, output o);
  assign o = i;
endmodule
