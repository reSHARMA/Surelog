module test (input size);
    logic [size:0][size-1:0] foo;
endmodule
